package yapp_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab7/Task1_data/sv/yapp_packet.sv"

endpackage